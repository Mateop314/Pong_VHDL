library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	
entity matrix_controller is 
end entity;

architecture rtl of matrix_controller is 
begin 

end architecture;